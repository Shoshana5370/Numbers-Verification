interface num_if(input logic clk,reset);
  
  logic [1:0] mytype;
  logic [15:0] data_in;
  logic [15:0] data_out;  
  
endinterface